module Jump_Controller(BranchE, func3, );


endmodule